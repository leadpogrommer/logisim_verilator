`ifndef CDM16_COMMON
`define CDM16_COMMON


localparam UC_ALU_ASRTD = 0;
localparam UC_DATA = 1;
localparam UC_FP_ASRT0 = 2;
localparam UC_IMM_ASRT1 = 3;
localparam UC_IMM_ASRTD = 4;
localparam UC_IMM_EXTEND_NEGATIVE = 5;
localparam UC_IMM_SHIFT = 6;
localparam UC_MEM = 7;
localparam UC_PC_ASRT0 = 8;
localparam UC_PC_ASRTD = 9;
localparam UC_PC_INC = 10;
localparam UC_PC_LATCH = 11;
localparam UC_PS_ASRTD = 12;
localparam UC_PS_LATCH_FLAGS = 13;
localparam UC_PS_LATCH_WORD = 14;
localparam UC_R_ASRT0 = 15;
localparam UC_R_ASRT1 = 16;
localparam UC_R_ASRTD = 17;
localparam UC_RLATCH = 18;
localparam UC_READ = 19;
localparam UC_SIGN_EXTEND = 20;
localparam UC_SP_ASRT0 = 21;
localparam UC_SP_ASRTD = 22;
localparam UC_SP_DEC = 23;
localparam UC_SP_INC = 24;
localparam UC_SP_LATCH = 25;
localparam UC_WORD = 26;
localparam UC_CUT = 27;

`endif