`timescale 1ns / 1ps


module color_bar(
    input                 clk,           //pixel clock
	input                 rst,           //reset signal high active
	output                hs,            //horizontal synchronization
	output                vs,            //vertical synchronization
	output                de,            //video valid
	output[7:0]           rgb_r,         //video red data
	output[7:0]           rgb_g,         //video green data
	output[7:0]           rgb_b,          //video blue data
	input [9:0]           char_line_data,
	output [12:0]         font_ram_addr,

    input [15:0] vram_data_in,
    output reg [15:0] vram_addr_in
);
 
//video timing parameter definition
//800x600 40Mhz
parameter H_ACTIVE = 16'd800; 
parameter H_FP = 16'd40;      
parameter H_SYNC = 16'd128;   
parameter H_BP = 16'd88;      
parameter V_ACTIVE = 16'd600; 
parameter V_FP  = 16'd1;     
parameter V_SYNC  = 16'd4;    
parameter V_BP  = 16'd23;    
parameter HS_POL = 1'b1;
parameter VS_POL = 1'b1;

 

parameter H_TOTAL = H_ACTIVE + H_FP + H_SYNC + H_BP;//horizontal total time (pixels)
parameter V_TOTAL = V_ACTIVE + V_FP + V_SYNC + V_BP;//vertical total time (lines)

reg hs_reg;                      //horizontal sync register
reg vs_reg;                      //vertical sync register
reg hs_reg_d0;                   //delay 1 clock of 'hs_reg'
reg vs_reg_d0;                   //delay 1 clock of 'vs_reg'
reg[11:0] h_cnt;                 //horizontal counter
reg[11:0] v_cnt;                 //vertical counter
reg[11:0] active_x;              //video x position 
reg[11:0] active_y;              //video y position 
reg[7:0] rgb_r_reg;              //video red data register
reg[7:0] rgb_g_reg;              //video green data register
reg[7:0] rgb_b_reg;              //video blue data register
reg h_active;                    //horizontal video active
reg v_active;                    //vertical video active
wire video_active;               //video active(horizontal active and vertical active)
reg video_active_d0;             //delay 1 clock of video_active
assign hs = hs_reg_d0;
assign vs = vs_reg_d0;
assign video_active = h_active & v_active;
assign de = video_active_d0;
assign rgb_r = rgb_r_reg;
assign rgb_g = rgb_g_reg;
assign rgb_b = rgb_b_reg;
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		begin
			hs_reg_d0 <= 1'b0;
			vs_reg_d0 <= 1'b0;
			video_active_d0 <= 1'b0;
		end
	else
		begin
			hs_reg_d0 <= hs_reg;
			vs_reg_d0 <= vs_reg;
			video_active_d0 <= video_active;
		end
end
 
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		h_cnt <= 12'd0;
	else if(h_cnt == H_TOTAL - 1)//horizontal counter maximum value
		h_cnt <= 12'd0;
	else
		h_cnt <= h_cnt + 12'd1;
end
 
 // char Width = 800/80 = 10
 // char Height = 600/30 = 20
 reg [6:0] char_x;
 reg [4:0] char_y;
 
 reg [4:0] char_pixel_line;
 reg [3:0] char_pixel_col;
 
 wire [7:0] char_num = char_y*80+char_x;
 
//  assign font_ram_addr = {char_num, char_pixel_line};
reg [16:0] char_data_latch;
reg [9:0] char_line_data_latch;

assign font_ram_addr = {vram_data_in[7:0], char_pixel_line};

// current x calculation
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		active_x <= 12'd0;
	else if(h_cnt >= H_FP + H_SYNC + H_BP - 1)//horizontal video active
		active_x <= h_cnt - (H_FP[11:0] + H_SYNC[11:0] + H_BP[11:0] - 12'd1);
	else
		active_x <= active_x;
	
	if(rst == 1'b1 || (h_cnt == H_FP + H_SYNC + H_BP - 1 - 10)) begin
	   char_x <= 127;
	   char_pixel_col <= 0;
	end else begin

        if (char_pixel_col == 1) begin
             char_x <= char_x + 1;
             vram_addr_in <= char_y*80+((char_x+1)&8'b01111111);
        end 

	   if(char_pixel_col == 9) begin
	       char_pixel_col <= 0;
           char_line_data_latch <= char_line_data;
           char_data_latch <= vram_data_in;
       end else begin
            char_pixel_col <= char_pixel_col + 1;
       end
	end
	
	
end
 
// current y calculation
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1) begin
		v_cnt <= 12'd0;
	    char_y = 0;
	    char_pixel_line = 0;
	end else if(h_cnt == H_FP  - 1)//horizontal sync time
		if(v_cnt == V_TOTAL - 1) begin//vertical counter maximum value
			v_cnt <= 12'd0;
			   
		end else begin
		    v_cnt <= v_cnt + 12'd1;
		    
		    if (v_cnt == V_FP + V_SYNC + V_BP - 1) begin
		       char_y = 0;
	           char_pixel_line = 0;
	         end else begin
                if (char_pixel_line == 19) begin
                  char_pixel_line <= 0;
                  char_y <= char_y + 1;
                end else char_pixel_line <= char_pixel_line + 1;
		    end
		end
	else
		v_cnt <= v_cnt;
end
 
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		hs_reg <= 1'b0;
	else if(h_cnt == H_FP - 1)//horizontal sync begin
		hs_reg <= HS_POL;
	else if(h_cnt == H_FP + H_SYNC - 1)//horizontal sync end
		hs_reg <= ~hs_reg;
	else
		hs_reg <= hs_reg;
end
 
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		h_active <= 1'b0;
	else if(h_cnt == H_FP + H_SYNC + H_BP - 1)//horizontal active begin
		h_active <= 1'b1;
	else if(h_cnt == H_TOTAL - 1)//horizontal active end
		h_active <= 1'b0;
	else
		h_active <= h_active;
end
 
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		vs_reg <= 1'd0;
	else if((v_cnt == V_FP - 1) && (h_cnt == H_FP - 1))//vertical sync begin
		vs_reg <= HS_POL;
	else if((v_cnt == V_FP + V_SYNC - 1) && (h_cnt == H_FP - 1))//vertical sync end
		vs_reg <= ~vs_reg;  
	else
		vs_reg <= vs_reg;
end
 
 reg [11:0] frame_cntr;
 
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		v_active <= 1'd0;
	else if((v_cnt == V_FP + V_SYNC + V_BP - 1) && (h_cnt == H_FP - 1))//vertical active begin
		begin 
		v_active <= 1'b1;
		frame_cntr <= frame_cntr + 1;
		end
	else if((v_cnt == V_TOTAL - 1) && (h_cnt == H_FP - 1)) //vertical active end
		v_active <= 1'b0;   
	else
		v_active <= v_active;
end

wire pixel_data = char_line_data_latch[char_pixel_col];
 
wire [7:0] char_style = char_data_latch[15:8];

wire is_dim = char_style[6];
wire is_blink = char_style[7];
wire [2:0] bg_color = char_style[5:3];
wire [2:0] fg_color = char_style[2:0];

wire [7:0] rgb_res [2:0];

genvar chan;
generate
    for(chan = 0; chan < 3; chan = chan + 1) begin
        assign rgb_res[chan] = {8{pixel_data ? (!fg_color[chan]) : (bg_color[chan])}} & {!is_dim, 7'b1111111} & {8{(!is_blink) | (frame_cntr[4])}};
    end
endgenerate
 
always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		begin
			rgb_r_reg <= 8'h00;
			rgb_g_reg <= 8'h00;
			rgb_b_reg <= 8'h00;
		end
	else if(video_active) begin	
            // TODO: I think these are messed up in hardware
          rgb_r_reg <= rgb_res[0];
          rgb_g_reg <= rgb_res[2];
          rgb_b_reg <= rgb_res[1];
	end else
		begin
			rgb_r_reg <= 8'h00;
			rgb_g_reg <= 8'h00;
			rgb_b_reg <= 8'h00;
		end
end
endmodule
